///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: Grounder
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();

reg myInput;

Grounder myGrounder(myInput);

initial begin
///////////////////////////////////////////////////////////////////////////////////
// Inputs: myInput (1 bit)
myInput=1; #10; 
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// No output to test
// Just really checking to make sure it doesn't crash
$display("All tests passed.");
///////////////////////////////////////////////////////////////////////////////////
end

endmodule
